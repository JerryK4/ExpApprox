library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity microprocessor is
    port (
        clk         : in  std_logic;
        rst         : in  std_logic;
        start       : in  std_logic;
        
        -- Giao ti?p v?i Unified Memory
        mem_data_in : in  std_logic_vector(15 downto 0); -- D? li?u ??c t? Memory (z_init)
        mem_addr    : out std_logic_vector(5 downto 0);  -- ??a ch? g?i t?i Memory
        mem_data_out: out std_logic_vector(15 downto 0); -- D? li?u ghi v�o Memory (exp_out)
        Mre         : out std_logic;
        Mwe         : out std_logic;
        
        done        : out std_logic
    );
end microprocessor;

architecture structural of microprocessor is

    --------------------------------------------------------------------
    -- COMPONENT DECLARATIONS
    --------------------------------------------------------------------
    component control_unit is
        port (
            clk      : in  std_logic;
            rst      : in  std_logic;
            start    : in  std_logic;
            rs       : in  std_logic;
            cal      : in  std_logic;

            x_sel    : out std_logic_vector(1 downto 0);
            y_sel    : out std_logic_vector(1 downto 0);
            z_sel    : out std_logic_vector(1 downto 0);
            i_sel    : out std_logic;
            x_en     : out std_logic;
            y_en     : out std_logic;
            z_en     : out std_logic;
            i_en     : out std_logic;

            Mre      : out std_logic;
            Mwe      : out std_logic;
            address  : out std_logic_vector(5 downto 0);
            done     : out std_logic
        );
    end component;

    component datapath is
        port(
            clk     : in std_logic;
            rst     : in std_logic;
            x_sel   : in std_logic_vector(1 downto 0);
            y_sel   : in std_logic_vector(1 downto 0);
            z_sel   : in std_logic_vector(1 downto 0);
            i_sel   : in std_logic;
            x_en    : in std_logic;
            y_en    : in std_logic;
            z_en    : in std_logic;
            i_en    : in std_logic;
            i_in    : in std_logic_vector(4 downto 0); 
            x_in    : in std_logic_vector(15 downto 0); 
            y_in    : in std_logic_vector(15 downto 0); 
            z_in    : in std_logic_vector(15 downto 0); 
            cal     : out std_logic;
            rs      : out std_logic;
            exp_out : out std_logic_vector(15 downto 0)
        );
    end component;

    --------------------------------------------------------------------
    -- INTERNAL SIGNALS (Control Signals & Status Flags)
    --------------------------------------------------------------------
    signal s_x_sel, s_y_sel, s_z_sel : std_logic_vector(1 downto 0);
    signal s_i_sel                   : std_logic;
    signal s_x_en, s_y_en, s_z_en    : std_logic;
    signal s_i_en	             : std_logic;
    signal s_rs, s_cal               : std_logic;

    -- CORDIC Constants (Q3.13)
    -- X_INIT = 1/Ke (H? s? t? l? Hyperbolic CORDIC)
    constant X_INIT_VAL : std_logic_vector(15 downto 0) := x"2690"; 
    constant Y_INIT_VAL : std_logic_vector(15 downto 0) := x"0000";
    constant I_START    : std_logic_vector(4 downto 0)  := "00001"; -- B?t ??u t? i=1

begin

    --------------------------------------------------------------------
    -- CONTROL UNIT INSTANTIATION
    --------------------------------------------------------------------
    U_CU: control_unit
        port map (
            clk      => clk,
            rst      => rst,
            start    => start,
            rs       => s_rs,
            cal      => s_cal,

            x_sel    => s_x_sel,
            y_sel    => s_y_sel,
            z_sel    => s_z_sel,
            i_sel    => s_i_sel,
            x_en     => s_x_en,
            y_en     => s_y_en,
            z_en     => s_z_en,
            i_en     => s_i_en,

            Mre      => Mre,
            Mwe      => Mwe,
            address  => mem_addr,
            done     => done
        );

    --------------------------------------------------------------------
    -- DATAPATH INSTANTIATION
    --------------------------------------------------------------------
    U_DP: datapath
        port map (
            clk     => clk,
            rst     => rst,
            
            x_sel   => s_x_sel,
            y_sel   => s_y_sel,
            z_sel   => s_z_sel,
            i_sel   => s_i_sel,
            
            x_en    => s_x_en,
            y_en    => s_y_en,
            z_en    => s_z_en,
            i_en    => s_i_en,

            i_in    => I_START,
            x_in    => X_INIT_VAL,
            y_in    => Y_INIT_VAL,
            z_in    => mem_data_in, -- L?y t? b? nh?

            cal     => s_cal,
            rs      => s_rs,
            exp_out => mem_data_out -- G?i k?t qu? v? b? nh?
        );

end structural;
